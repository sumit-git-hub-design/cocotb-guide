`timescale 1ns/1ps

module mux();

endmodule
