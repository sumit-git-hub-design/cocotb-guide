`timescale 1ns/1ps

module mux();

initial begin
  $display("This display is present in DUT");
end

endmodule
